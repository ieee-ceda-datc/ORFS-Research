# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0050 ;

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER active
  TYPE MASTERSLICE ;
END active

LAYER M1
  TYPE ROUTING ;
  SPACING 0.065 ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  HEIGHT 0.37 ;
  CAPACITANCE CPERSQDIST 7.7161e-05 ;
  EDGECAPACITANCE 2.7365e-05 ;
END M1

LAYER via1
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via1

LAYER M2
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.62 ;
  CAPACITANCE CPERSQDIST 4.0896e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M2

LAYER via2
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via2

LAYER M3
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M3

LAYER via3
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via3

LAYER M4
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.14 ;
  CAPACITANCE CPERSQDIST 2.0743e-05 ;
  EDGECAPACITANCE 3.0908e-05 ;
END M4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via4

LAYER M5
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.71 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 2.3863e-06 ;
END M5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via5

LAYER M6
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 2.28 ;
  CAPACITANCE CPERSQDIST 1.0036e-05 ;
  EDGECAPACITANCE 2.3863e-05 ;
END M6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via6

LAYER M7
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 2.85 ;
  CAPACITANCE CPERSQDIST 7.9771e-06 ;
  EDGECAPACITANCE 3.2577e-05 ;
END M7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via7

LAYER M8
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 4.47 ;
  CAPACITANCE CPERSQDIST 5.0391e-06 ;
  EDGECAPACITANCE 2.3932e-05 ;
END M8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via8

LAYER M9
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 6.09 ;
  CAPACITANCE CPERSQDIST 3.6827e-06 ;
  EDGECAPACITANCE 3.0803e-05 ;
END M9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  RESISTANCE 0.5 ;
END via9

LAYER M10
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 10.09 ;
  CAPACITANCE CPERSQDIST 2.2124e-06 ;
  EDGECAPACITANCE 2.3667e-05 ;
END M10

LAYER hb_layer
  TYPE CUT ;
  SPACING 1.8 ;
  WIDTH 1.2 ;
  RESISTANCE 0.02 ;
END hb_layer

LAYER M12
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 6.09 ;
  CAPACITANCE CPERSQDIST 3.6827e-06 ;
  EDGECAPACITANCE 3.0803e-05 ;
END M12

LAYER via12
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via12

LAYER M13
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 4.47 ;
  CAPACITANCE CPERSQDIST 5.0391e-06 ;
  EDGECAPACITANCE 2.3932e-05 ;
END M13

LAYER via13
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via13

LAYER M14
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 2.85 ;
  CAPACITANCE CPERSQDIST 7.9771e-06 ;
  EDGECAPACITANCE 3.2577e-05 ;
END M14

LAYER via14
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via14

LAYER M15
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 2.28 ;
  CAPACITANCE CPERSQDIST 1.0036e-05 ;
  EDGECAPACITANCE 2.3863e-05 ;
END M15

LAYER via15
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via15

LAYER M16
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.71 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 2.3863e-06 ;
END M16

LAYER via16
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via16

LAYER M17
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.14 ;
  CAPACITANCE CPERSQDIST 2.0743e-05 ;
  EDGECAPACITANCE 3.0908e-05 ;
END M17

LAYER via17
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via17

LAYER M18
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M18

LAYER via18
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via18

LAYER M19
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.62 ;
  CAPACITANCE CPERSQDIST 4.0896e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M19

LAYER via19
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via19

LAYER M20
  TYPE ROUTING ;
  SPACING 0.065 ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  HEIGHT 0.37 ;
  CAPACITANCE CPERSQDIST 7.7161e-05 ;
  EDGECAPACITANCE 2.7365e-05 ;
END M20

LAYER via20
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via20

LAYER M21
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.62 ;
  CAPACITANCE CPERSQDIST 4.0896e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M21

LAYER via21
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via21

LAYER M22
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M22

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA via1_4 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_4

VIA via1_0 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_0

VIA via1_1 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_1

VIA via1_2 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_2

VIA via1_3 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_3

VIA via1_5 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_5

VIA via1_6 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_6

VIA via1_7 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_7

VIA via1_8 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_8

VIA via2_8 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_8

VIA via2_4 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_4

VIA via2_5 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_5

VIA via2_7 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_7

VIA via2_6 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_6

VIA via2_0 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_0

VIA via2_1 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_1

VIA via2_2 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_2

VIA via2_3 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_3

VIA via3_2 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_2

VIA via3_0 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_0

VIA via3_1 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_1

VIA via4_0 DEFAULT
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4_0

VIA via5_0 DEFAULT
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5_0

VIA via6_0 DEFAULT
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via6_0

VIA via7_0 DEFAULT
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via7_0

VIA via8_0 DEFAULT
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via8_0

VIA via9_0 DEFAULT
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via9_0

VIA hb_layer_0 DEFAULT
  LAYER hb_layer ;
    RECT -0.6 -0.6 0.6 0.6 ;
  LAYER M10 ;
    RECT -0.6 -0.6 0.6 0.6 ;
  LAYER M12 ;
    RECT -0.6 -0.6 0.6 0.6 ;
END hb_layer_0

VIA via12_0 DEFAULT
  LAYER via12 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M12 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M13 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via12_0

VIA via13_0 DEFAULT
  LAYER via13 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M13 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M14 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via13_0

VIA via14_0 DEFAULT
  LAYER via14 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M14 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M15 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via14_0

VIA via15_0 DEFAULT
  LAYER via15 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M15 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M16 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via15_0

VIA via16_0 DEFAULT
  LAYER via16 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M16 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M17 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via16_0

VIA via17_2 DEFAULT
  LAYER via17 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M17 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via17_2

VIA via17_0 DEFAULT
  LAYER via17 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M17 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M18 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via17_0

VIA via17_1 DEFAULT
  LAYER via17 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M17 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M18 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via17_1

VIA via18_8 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via18_8

VIA via18_4 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M19 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via18_4

VIA via18_5 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M19 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via18_5

VIA via18_7 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M19 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via18_7

VIA via18_6 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via18_6

VIA via18_0 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M19 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via18_0

VIA via18_1 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M19 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via18_1

VIA via18_2 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M19 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via18_2

VIA via18_3 DEFAULT
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M18 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M19 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via18_3

VIA via19_4 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M20 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via19_4

VIA via19_0 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M20 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via19_0

VIA via19_1 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M20 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via19_1

VIA via19_2 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M20 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via19_2

VIA via19_3 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M20 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via19_3

VIA via19_5 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M20 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via19_5

VIA via19_6 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via19_6

VIA via19_7 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M20 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via19_7

VIA via19_8 DEFAULT
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M19 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via19_8

VIA via20_4 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M21 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via20_4

VIA via20_0 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M21 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via20_0

VIA via20_1 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M21 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via20_1

VIA via20_2 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M21 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via20_2

VIA via20_3 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M21 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via20_3

VIA via20_5 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M21 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via20_5

VIA via20_6 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via20_6

VIA via20_7 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M21 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via20_7

VIA via20_8 DEFAULT
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M20 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via20_8

VIA via21_8 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M22 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via21_8

VIA via21_4 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M22 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via21_4

VIA via21_5 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M22 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via21_5

VIA via21_7 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M22 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via21_7

VIA via21_6 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via21_6

VIA via21_0 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via21_0

VIA via21_1 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M22 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via21_1

VIA via21_2 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M22 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via21_2

VIA via21_3 DEFAULT
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M21 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via21_3

VIARULE Via1Array-0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-0

VIARULE Via1Array-1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-1

VIARULE Via1Array-2 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-2

VIARULE Via1Array-3 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-3

VIARULE Via1Array-4 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0 ;
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-4

VIARULE Via2Array-0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-0

VIARULE Via2Array-1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-1

VIARULE Via2Array-2 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-2

VIARULE Via2Array-3 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-3

VIARULE Via2Array-4 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER M3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-4

VIARULE Via3Array-0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-0

VIARULE Via3Array-1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.035 ;
  LAYER M4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-1

VIARULE Via3Array-2 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.035 0 ;
  LAYER M4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-2

VIARULE Via4Array-0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0 ;
  LAYER M5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-0

VIARULE Via5Array-0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0 0 ;
  LAYER M6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-0

VIARULE Via6Array-0 GENERATE
  LAYER M6 ;
    ENCLOSURE 0 0 ;
  LAYER M7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-0

VIARULE Via7Array-0 GENERATE
  LAYER M7 ;
    ENCLOSURE 0 0 ;
  LAYER M8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-0

VIARULE Via8Array-0 GENERATE
  LAYER M8 ;
    ENCLOSURE 0 0 ;
  LAYER M9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-0

VIARULE Via9Array-0 GENERATE
  LAYER M10 ;
    ENCLOSURE 0 0 ;
  LAYER M9 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-0

VIARULE hb_layerArray-0 GENERATE
  LAYER M12 ;
    ENCLOSURE 0 0 ;
  LAYER M10 ;
    ENCLOSURE 0 0 ;
  LAYER hb_layer ;
    RECT -0.6 -0.6 0.6 0.6 ;
    SPACING 3.0 BY 3.0 ;
END hb_layerArray-0

VIARULE Via12Array-0 GENERATE
  LAYER M12 ;
    ENCLOSURE 0 0 ;
  LAYER M13 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via12 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via12Array-0

VIARULE Via13Array-0 GENERATE
  LAYER M13 ;
    ENCLOSURE 0 0 ;
  LAYER M14 ;
    ENCLOSURE 0 0 ;
  LAYER via13 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via13Array-0

VIARULE Via14Array-0 GENERATE
  LAYER M14 ;
    ENCLOSURE 0 0 ;
  LAYER M15 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via14 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via14Array-0

VIARULE Via15Array-0 GENERATE
  LAYER M15 ;
    ENCLOSURE 0 0 ;
  LAYER M16 ;
    ENCLOSURE 0 0 ;
  LAYER via15 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via15Array-0

VIARULE Via16Array-0 GENERATE
  LAYER M16 ;
    ENCLOSURE 0 0 ;
  LAYER M17 ;
    ENCLOSURE 0 0 ;
  LAYER via16 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via16Array-0

VIARULE Via17Array-0 GENERATE
  LAYER M17 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M18 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via17 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via17Array-0

VIARULE Via17Array-1 GENERATE
  LAYER M17 ;
    ENCLOSURE 0 0.035 ;
  LAYER M18 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via17 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via17Array-1

VIARULE Via17Array-2 GENERATE
  LAYER M17 ;
    ENCLOSURE 0.035 0 ;
  LAYER M18 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via17 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via17Array-2

VIARULE Via18Array-0 GENERATE
  LAYER M18 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M19 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via18Array-0

VIARULE Via18Array-1 GENERATE
  LAYER M18 ;
    ENCLOSURE 0 0.035 ;
  LAYER M19 ;
    ENCLOSURE 0 0.035 ;
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via18Array-1

VIARULE Via18Array-2 GENERATE
  LAYER M18 ;
    ENCLOSURE 0.035 0 ;
  LAYER M19 ;
    ENCLOSURE 0.035 0 ;
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via18Array-2

VIARULE Via18Array-3 GENERATE
  LAYER M18 ;
    ENCLOSURE 0 0.035 ;
  LAYER M19 ;
    ENCLOSURE 0.035 0 ;
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via18Array-3

VIARULE Via18Array-4 GENERATE
  LAYER M18 ;
    ENCLOSURE 0.035 0 ;
  LAYER M19 ;
    ENCLOSURE 0 0.035 ;
  LAYER via18 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via18Array-4

VIARULE Via19Array-0 GENERATE
  LAYER M19 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M20 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via19Array-0

VIARULE Via19Array-1 GENERATE
  LAYER M19 ;
    ENCLOSURE 0 0.035 ;
  LAYER M20 ;
    ENCLOSURE 0 0.035 ;
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via19Array-1

VIARULE Via19Array-2 GENERATE
  LAYER M19 ;
    ENCLOSURE 0.035 0 ;
  LAYER M20 ;
    ENCLOSURE 0.035 0 ;
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via19Array-2

VIARULE Via19Array-3 GENERATE
  LAYER M19 ;
    ENCLOSURE 0 0.035 ;
  LAYER M20 ;
    ENCLOSURE 0.035 0 ;
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via19Array-3

VIARULE Via19Array-4 GENERATE
  LAYER M19 ;
    ENCLOSURE 0.035 0 ;
  LAYER M20 ;
    ENCLOSURE 0 0.035 ;
  LAYER via19 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via19Array-4

VIARULE Via20Array-0 GENERATE
  LAYER M20 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M21 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via20Array-0

VIARULE Via20Array-1 GENERATE
  LAYER M20 ;
    ENCLOSURE 0 0.035 ;
  LAYER M21 ;
    ENCLOSURE 0 0.035 ;
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via20Array-1

VIARULE Via20Array-2 GENERATE
  LAYER M20 ;
    ENCLOSURE 0.035 0 ;
  LAYER M21 ;
    ENCLOSURE 0.035 0 ;
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via20Array-2

VIARULE Via20Array-3 GENERATE
  LAYER M20 ;
    ENCLOSURE 0 0.035 ;
  LAYER M21 ;
    ENCLOSURE 0.035 0 ;
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via20Array-3

VIARULE Via20Array-4 GENERATE
  LAYER M20 ;
    ENCLOSURE 0.035 0 ;
  LAYER M21 ;
    ENCLOSURE 0 0.035 ;
  LAYER via20 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via20Array-4

VIARULE Via21Array-0 GENERATE
  LAYER M21 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M22 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via21Array-0

VIARULE Via21Array-1 GENERATE
  LAYER M21 ;
    ENCLOSURE 0 0.035 ;
  LAYER M22 ;
    ENCLOSURE 0 0.035 ;
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via21Array-1

VIARULE Via21Array-2 GENERATE
  LAYER M21 ;
    ENCLOSURE 0.035 0 ;
  LAYER M22 ;
    ENCLOSURE 0.035 0 ;
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via21Array-2

VIARULE Via21Array-3 GENERATE
  LAYER M21 ;
    ENCLOSURE 0 0.035 ;
  LAYER M22 ;
    ENCLOSURE 0.035 0 ;
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via21Array-3

VIARULE Via21Array-4 GENERATE
  LAYER M21 ;
    ENCLOSURE 0.035 0 ;
  LAYER M22 ;
    ENCLOSURE 0 0.035 ;
  LAYER via21 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via21Array-4

SPACING
  SAMENET M1 M1 0.065 ;
  SAMENET M2 M2 0.07 ;
  SAMENET M3 M3 0.07 ;
  SAMENET M4 M4 0.14 ;
  SAMENET M5 M5 0.14 ;
  SAMENET M6 M6 0.14 ;
  SAMENET M7 M7 0.4 ;
  SAMENET M8 M8 0.4 ;
  SAMENET M9 M9 0.8 ;
  SAMENET M10 M10 0.8 ;
  SAMENET M12 M12 0.8 ;
  SAMENET M13 M13 0.4 ;
  SAMENET M14 M14 0.4 ;
  SAMENET M15 M15 0.14 ;
  SAMENET M16 M16 0.14 ;
  SAMENET M17 M17 0.14 ;
  SAMENET M18 M18 0.07 ;
  SAMENET M19 M19 0.07 ;
  SAMENET M20 M20 0.065 ;
  SAMENET M21 M21 0.07 ;
  SAMENET M22 M22 0.07 ;
  SAMENET via1 via1 0.08 ;
  SAMENET via2 via2 0.09 ;
  SAMENET via3 via3 0.09 ;
  SAMENET via4 via4 0.16 ;
  SAMENET via5 via5 0.16 ;
  SAMENET via6 via6 0.16 ;
  SAMENET via7 via7 0.44 ;
  SAMENET via8 via8 0.44 ;
  SAMENET via9 via9 0.88 ;
  SAMENET hb_layer hb_layer 1.8 ;
  SAMENET via12 via12 0.44 ;
  SAMENET via13 via13 0.44 ;
  SAMENET via14 via14 0.16 ;
  SAMENET via15 via15 0.16 ;
  SAMENET via16 via16 0.16 ;
  SAMENET via17 via17 0.09 ;
  SAMENET via18 via18 0.09 ;
  SAMENET via19 via19 0.08 ;
  SAMENET via20 via20 0.08 ;
  SAMENET via21 via21 0.09 ;
  SAMENET via1 via2 0.0 STACK ;
  SAMENET via2 via3 0.0 STACK ;
  SAMENET via3 via4 0.0 STACK ;
  SAMENET via4 via5 0.0 STACK ;
  SAMENET via5 via6 0.0 STACK ;
  SAMENET via6 via7 0.0 STACK ;
  SAMENET via7 via8 0.0 STACK ;
  SAMENET via8 via9 0.0 STACK ;
  SAMENET via9 hb_layer 0.0 STACK ;
  SAMENET hb_layer via12 0.0 STACK ;
  SAMENET via12 via13 0.0 STACK ;
  SAMENET via13 via14 0.0 STACK ;
  SAMENET via14 via15 0.0 STACK ;
  SAMENET via15 via16 0.0 STACK ;
  SAMENET via16 via17 0.0 STACK ;
  SAMENET via17 via18 0.0 STACK ;
  SAMENET via18 via19 0.0 STACK ;
  SAMENET via19 via20 0.0 STACK ;
  SAMENET via20 via21 0.0 STACK ;
END SPACING

SITE FreePDK45_38x28_10R_NP_162NW_34O
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 1.4 ;
END FreePDK45_38x28_10R_NP_162NW_34O

END LIBRARY
#
# End of file
#
