VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x15_upper
  FOREIGN fakeram45_64x15_upper 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 11.210 BY 58.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 12.880 0.070 12.950 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 14.560 0.070 14.630 ;
    END
  END w_mask_in[14]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 16.240 0.070 16.310 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 17.920 0.070 17.990 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 19.600 0.070 19.670 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 20.440 0.070 20.510 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 21.280 0.070 21.350 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 22.120 0.070 22.190 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END rd_out[14]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 29.680 0.070 29.750 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 30.520 0.070 30.590 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 31.360 0.070 31.430 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 33.040 0.070 33.110 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 34.720 0.070 34.790 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 36.400 0.070 36.470 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 37.240 0.070 37.310 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 38.080 0.070 38.150 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 38.920 0.070 38.990 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 39.760 0.070 39.830 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 40.600 0.070 40.670 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 41.440 0.070 41.510 ;
    END
  END wd_in[14]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 43.120 0.070 43.190 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 43.960 0.070 44.030 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 44.800 0.070 44.870 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 45.640 0.070 45.710 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 46.480 0.070 46.550 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 47.320 0.070 47.390 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 49.840 0.070 49.910 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 50.680 0.070 50.750 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M17 ;
      RECT 2.660 2.800 2.940 56.000 ;
      RECT 7.140 2.800 7.420 56.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M17 ;
      RECT 4.900 2.800 5.180 56.000 ;
    END
  END VDD
  OBS
    LAYER M20 ;
    RECT 0 0 11.210 58.800 ;
    LAYER M19 ;
    RECT 0 0 11.210 58.800 ;
    LAYER M18 ;
    RECT 0.070 0 11.210 58.800 ;
    RECT 0 0.000 0.070 2.800 ;
    RECT 0 2.870 0.070 3.640 ;
    RECT 0 3.710 0.070 4.480 ;
    RECT 0 4.550 0.070 5.320 ;
    RECT 0 5.390 0.070 6.160 ;
    RECT 0 6.230 0.070 7.000 ;
    RECT 0 7.070 0.070 7.840 ;
    RECT 0 7.910 0.070 8.680 ;
    RECT 0 8.750 0.070 9.520 ;
    RECT 0 9.590 0.070 10.360 ;
    RECT 0 10.430 0.070 11.200 ;
    RECT 0 11.270 0.070 12.040 ;
    RECT 0 12.110 0.070 12.880 ;
    RECT 0 12.950 0.070 13.720 ;
    RECT 0 13.790 0.070 14.560 ;
    RECT 0 14.630 0.070 16.240 ;
    RECT 0 16.310 0.070 17.080 ;
    RECT 0 17.150 0.070 17.920 ;
    RECT 0 17.990 0.070 18.760 ;
    RECT 0 18.830 0.070 19.600 ;
    RECT 0 19.670 0.070 20.440 ;
    RECT 0 20.510 0.070 21.280 ;
    RECT 0 21.350 0.070 22.120 ;
    RECT 0 22.190 0.070 22.960 ;
    RECT 0 23.030 0.070 23.800 ;
    RECT 0 23.870 0.070 24.640 ;
    RECT 0 24.710 0.070 25.480 ;
    RECT 0 25.550 0.070 26.320 ;
    RECT 0 26.390 0.070 27.160 ;
    RECT 0 27.230 0.070 28.000 ;
    RECT 0 28.070 0.070 29.680 ;
    RECT 0 29.750 0.070 30.520 ;
    RECT 0 30.590 0.070 31.360 ;
    RECT 0 31.430 0.070 32.200 ;
    RECT 0 32.270 0.070 33.040 ;
    RECT 0 33.110 0.070 33.880 ;
    RECT 0 33.950 0.070 34.720 ;
    RECT 0 34.790 0.070 35.560 ;
    RECT 0 35.630 0.070 36.400 ;
    RECT 0 36.470 0.070 37.240 ;
    RECT 0 37.310 0.070 38.080 ;
    RECT 0 38.150 0.070 38.920 ;
    RECT 0 38.990 0.070 39.760 ;
    RECT 0 39.830 0.070 40.600 ;
    RECT 0 40.670 0.070 41.440 ;
    RECT 0 41.510 0.070 43.120 ;
    RECT 0 43.190 0.070 43.960 ;
    RECT 0 44.030 0.070 44.800 ;
    RECT 0 44.870 0.070 45.640 ;
    RECT 0 45.710 0.070 46.480 ;
    RECT 0 46.550 0.070 47.320 ;
    RECT 0 47.390 0.070 49.000 ;
    RECT 0 49.070 0.070 49.840 ;
    RECT 0 49.910 0.070 50.680 ;
    RECT 0 50.750 0.070 58.800 ;
    LAYER M17 ;
    RECT 0 0 11.210 2.800 ;
    RECT 0 56.000 11.210 58.800 ;
    RECT 0.000 2.800 2.660 56.000 ;
    RECT 2.940 2.800 4.900 56.000 ;
    RECT 5.180 2.800 7.140 56.000 ;
    RECT 7.420 2.800 11.210 56.000 ;
  END
END fakeram45_64x15_upper

END LIBRARY
